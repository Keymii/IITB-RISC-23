library std;
library ieee;
use std.standard.all;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity subCircuit_RR is
  port ( instr: in std_logic_vector(15 downto 0);

			reg_read_1: in STD_LOGIC;
			reg_read_2: in STD_LOGIC;
			
			rf_a1,rf_a2:out std_logic_vector(2 downto 0);
			rf_d1,rf_d2:in std_logic_vector(15 downto 0);
		 
    );
	 
end subCircuit_RR;
architecture a3 of subCircuit_RR is

begin

end a3;
 
 

 