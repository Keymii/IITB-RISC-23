library std;
library ieee;
use std.standard.all;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity subCircuit_EX is
  port ( instr: in std_logic_vector(15 downto 0);
				
		 
    );
	 
end subCircuit_EX;
architecture behav of subCircuit_EX is

begin

end behav;